// TITLE: convert_to_binary.sv
// PROJECT: Keyboard VLSI lab
// DESCRIPTION: Look-up-table

`timescale 1ns/1ps

module convert_to_binary (
    input logic [7:0] scan_code_in,
    output logic [3:0] binary_out
    );
    // Simple combinational logic using case statements (LUT)
endmodule
