// TITLE: binary_to_sgd.sv
// PROJECT: Keyboard VLSI lab
// DESCRIPTION: Simple look-up table

`timescale 1ns/1ps

module binary_to_sg (
    input logic [3:0] binary_in,
    output logic [7:0] sev_seg
    );

endmodule
